// lib for graphwiz
// to define input and outputs

module DL000D_4x1NAND2(output Y, input A, B);
endmodule

module DL002D_4x1NOR2(output Y, input A, B);
endmodule

module DL004D_6x1NOT(output Y, input A);
endmodule

module DL011D_3x1AND3(output Y, input A, B, C);
endmodule

module DL020D_2x1NAND4(output Y, input A, B, C, D);
endmodule

module DL032D_4x1OR2(output Y, input A, B);
endmodule

module DL086D_4x1XOR2(output Y, input A, B);
endmodule

module DL374D_8x1DFF(output Q, input CLK, D);
endmodule
